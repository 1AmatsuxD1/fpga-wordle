--------------------------------------------------------------------------------
-- Character ROM: เก็บ Bitmap Font สำหรับตัวอักษร A-Z
-- ขนาดตัวอักษร: 8×8 pixels ต่อตัว
-- รองรับ: A-Z (uppercase)
-- Clock: 20 MHz
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity char_rom is
    Port (
        clk       : in  std_logic;
        char_code : in  std_logic_vector(7 downto 0);  -- ASCII code (0x41-0x5A = A-Z)
        row       : in  unsigned(2 downto 0);          -- แถวที่ 0-7
        col       : in  unsigned(2 downto 0);          -- คอลัมน์ที่ 0-7
        pixel     : out std_logic                      -- 0=ไม่วาด, 1=วาด
    );
end char_rom;

architecture Behavioral of char_rom is
    
    -- ประเภทข้อมูล: แต่ละตัวอักษร = 8 แถว × 8 บิต
    type char_row is array (0 to 7) of std_logic_vector(7 downto 0);
    type font_rom is array (0 to 25) of char_row;
    
    -- Font ROM: 26 ตัวอักษร (A-Z)
    -- 1 = วาดพิกเซล, 0 = ไม่วาด
    constant FONT : font_rom := (
        -- A (index 0)
        0 => (
            x"18",  -- 00011000
            x"24",  -- 00100100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"7E",  -- 01111110
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"00"   -- 00000000
        ),
        
        -- B (index 1)
        1 => (
            x"7C",  -- 01111100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"7C",  -- 01111100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"7C",  -- 01111100
            x"00"   -- 00000000
        ),
        
        -- C (index 2)
        2 => (
            x"3C",  -- 00111100
            x"42",  -- 01000010
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"42",  -- 01000010
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- D (index 3)
        3 => (
            x"78",  -- 01111000
            x"44",  -- 01000100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"44",  -- 01000100
            x"78",  -- 01111000
            x"00"   -- 00000000
        ),
        
        -- E (index 4)
        4 => (
            x"7E",  -- 01111110
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"7C",  -- 01111100
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"7E",  -- 01111110
            x"00"   -- 00000000
        ),
        
        -- F (index 5)
        5 => (
            x"7E",  -- 01111110
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"7C",  -- 01111100
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"00"   -- 00000000
        ),
        
        -- G (index 6)
        6 => (
            x"3C",  -- 00111100
            x"42",  -- 01000010
            x"40",  -- 01000000
            x"4E",  -- 01001110
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- H (index 7)
        7 => (
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"7E",  -- 01111110
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"00"   -- 00000000
        ),
        
        -- I (index 8)
        8 => (
            x"3C",  -- 00111100
            x"18",  -- 00011000
            x"18",  -- 00011000
            x"18",  -- 00011000
            x"18",  -- 00011000
            x"18",  -- 00011000
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- J (index 9)
        9 => (
            x"1E",  -- 00011110
            x"0C",  -- 00001100
            x"0C",  -- 00001100
            x"0C",  -- 00001100
            x"0C",  -- 00001100
            x"4C",  -- 01001100
            x"38",  -- 00111000
            x"00"   -- 00000000
        ),
        
        -- K (index 10)
        10 => (
            x"44",  -- 01000100
            x"48",  -- 01001000
            x"50",  -- 01010000
            x"60",  -- 01100000
            x"50",  -- 01010000
            x"48",  -- 01001000
            x"44",  -- 01000100
            x"00"   -- 00000000
        ),
        
        -- L (index 11)
        11 => (
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"7E",  -- 01111110
            x"00"   -- 00000000
        ),
        
        -- M (index 12)
        12 => (
            x"42",  -- 01000010
            x"66",  -- 01100110
            x"5A",  -- 01011010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"00"   -- 00000000
        ),
        
        -- N (index 13)
        13 => (
            x"42",  -- 01000010
            x"62",  -- 01100010
            x"52",  -- 01010010
            x"4A",  -- 01001010
            x"46",  -- 01000110
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"00"   -- 00000000
        ),
        
        -- O (index 14)
        14 => (
            x"3C",  -- 00111100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- P (index 15)
        15 => (
            x"7C",  -- 01111100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"7C",  -- 01111100
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"40",  -- 01000000
            x"00"   -- 00000000
        ),
        
        -- Q (index 16)
        16 => (
            x"3C",  -- 00111100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"52",  -- 01010010
            x"4A",  -- 01001010
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- R (index 17)
        17 => (
            x"7C",  -- 01111100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"7C",  -- 01111100
            x"50",  -- 01010000
            x"48",  -- 01001000
            x"44",  -- 01000100
            x"00"   -- 00000000
        ),
        
        -- S (index 18)
        18 => (
            x"3C",  -- 00111100
            x"42",  -- 01000010
            x"40",  -- 01000000
            x"3C",  -- 00111100
            x"02",  -- 00000010
            x"42",  -- 01000010
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- T (index 19)
        19 => (
            x"FE",  -- 11111110
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"00"   -- 00000000
        ),
        
        -- U (index 20)
        20 => (
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"3C",  -- 00111100
            x"00"   -- 00000000
        ),
        
        -- V (index 21)
        21 => (
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"24",  -- 00100100
            x"18",  -- 00011000
            x"00"   -- 00000000
        ),
        
        -- W (index 22)
        22 => (
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"5A",  -- 01011010
            x"66",  -- 01100110
            x"42",  -- 01000010
            x"00"   -- 00000000
        ),
        
        -- X (index 23)
        23 => (
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"24",  -- 00100100
            x"18",  -- 00011000
            x"24",  -- 00100100
            x"42",  -- 01000010
            x"42",  -- 01000010
            x"00"   -- 00000000
        ),
        
        -- Y (index 24)
        24 => (
            x"82",  -- 10000010
            x"44",  -- 01000100
            x"28",  -- 00101000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"10",  -- 00010000
            x"00"   -- 00000000
        ),
        
        -- Z (index 25)
        25 => (
            x"7E",  -- 01111110
            x"02",  -- 00000010
            x"04",  -- 00000100
            x"18",  -- 00011000
            x"20",  -- 00100000
            x"40",  -- 01000000
            x"7E",  -- 01111110
            x"00"   -- 00000000
        )
    );
    
    signal char_index : integer range 0 to 25;
    signal char_data  : std_logic_vector(7 downto 0);
    
begin
    
    -- แปลง ASCII code เป็น index (A=0, B=1, ..., Z=25)
    process(char_code)
    begin
        if unsigned(char_code) >= x"41" and unsigned(char_code) <= x"5A" then
            -- Uppercase A-Z
            char_index <= to_integer(unsigned(char_code) - x"41");
        elsif unsigned(char_code) >= x"61" and unsigned(char_code) <= x"7A" then
            -- Lowercase a-z (แปลงเป็น uppercase)
            char_index <= to_integer(unsigned(char_code) - x"61");
        else
            -- ไม่ใช่ตัวอักษร = แสดงช่องว่าง
            char_index <= 0;
        end if;
    end process;
    
    -- อ่านข้อมูลจาก ROM
    process(clk)
    begin
        if rising_edge(clk) then
            -- อ่านแถวของตัวอักษร
            char_data <= FONT(char_index)(to_integer(row));
            
            -- อ่านบิตเฉพาะคอลัมน์
            pixel <= char_data(7 - to_integer(col));
        end if;
    end process;
    
end Behavioral;